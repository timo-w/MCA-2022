BZh91AY&SY��0 7߀Ryg����������` (�    4Tdh# ���  4��I�i�    @@ q�&�#F	���h�#@1�L��M`&i�L� �2hb14`��@	��24I�h�2	��	�&���M#aM�驀���x$�eЌ	&�$�X����:zY�$`�:���ګ�?�j�J~���}[^����_�^9���p~Ť�[����R�%�$���k�����u��E8->���dT5T���nj�
>��������p�j٧�=/���i>Y�v2ɖ�/�+.Z��d��=����d����,�����>-��ֵ�YծU{S���L�:mg���j��/k�����[�ٷwOӺ�g+�}��}�2�#>k����r��m���kƫ֝n���^�԰�A3�s�Hrj�'�u� %A�`��ח��P��7D�Խ8P轙kd�b����uE^����M�0���Q�CuQ�x�kU�e�iUd֊dY3|Ŵ�Y�
���𘛢�*j^���Z����9�4b���9�4]�4���=�/c��=��u���V,�U�UUUUUU�eԴh�<��:��2�ʙ�J�U�1j��V���n����f�>z̧�~��K�--2����tb��W)fm�Ce#���5\m��F�Hԡ�[uU�'*���,(�)@��0�P\Yg����cd6W�8B�F레�c�������U_�PJ�7�]�� p�3�!2��RX/<��ͦ�r���/&����Uil�~�[3��ss&�1,:��N8���5S�6��=e*�4��?�D�"z�{�?!R��q�ۛ���w8>t�:��2>d��Յ~s��l�iw;�[ߪ����RO��^^�=?�7:�<��)^�A�дe+�n�m�Y���m��Ds6w�Z�K�]�b�J)����LE�2d��ɲ^��F���S�nq����p���[�<xw˽/+4Ւ�]����Qb��9"��؊�XYii��m�K���73)�՜�|���~�1���gKt���+�y\tt�4_wQ����uT�1dk�¾�3�����ԪJsɓ6o�{L������6|󸧶&�i�{�?�o�Fնy��r���J�tgj7��JT��/1���R��fQy߯�8gU���ľ$�*Έ����g�����V��OK)�2���v��xZ˯9���3ԯ/A������PѴ�Q�*}�c�r�m��j�d)<��Z�aX�BYO/i�S,z�N▴�YM$�sdOŴhz�݆�6D����f������(��)R�).K�#�,J��tNM�%��K�3��ud�j���mV0��U/R�X�*vJ�ݬ�7��4V�b�IE�F�D��~(hi�4iFZ��kJ�G���<>�d+��J�3v%�}��Fs�T<W�,�9�g�c�'�>Ë�����&�YI���99#���˂�ȴQ��vέ{G�֋�;��I�pk�ʪ�?�t}O#��tq�:?z�:Y>aID��`QH��C�?y��ӣk��So����s���՜52l&�J�ȕ
���k�fKҳ����x]N���ӿ&M��y'f�߈�e3���*�+v���^�'Q���Q��3��b�NY���GC�M��6�h��m߭�x��Շ&�塔Mx�L���R7>���P�2Q�ѿ��&�-�$�6(�2�o3��C���pgZ�&S���05�l�������Q�n��O׳���Je�*��)Hx�zb7��]��BB�7\�