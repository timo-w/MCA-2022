BZh91AY&SY�F�q \_�Ryg����������`  �     !$�4�dLF�4   �C c��41�0�L �F��2d��bh�#0�0Mdh��� h�!� h2�  8ɓC�� �� �M4i��*H�A�6�L�hѨ�(i�৵OML��ʓS�(�D`$��ɂO�?WԺ:��h&���K�z����=U�S��O[�٫��3�O�nYx�]8�r�r�� �j�����I�V��Rl��5E8�?�F�uR1)*tP��n48�W������8;�3�ОG�^�����1Ŏ�/�6^-i�l�������b͵��Yj)���p�^_�Z֖um�^���3�V��nʘ2U��Y�������N�7ur�{�&Qƺz/��?�+f\�X0����>�p$N�ۖ�Zޑط�w�?��~ޮD��Z����x�#��Ȝ�T��>>�/�iP��oM��S
^���{1�lR�8ڗ�ĵx�E���}3ƕI���Z�#J�?�N+���q�z��Z�&�ȴі��x=f���}����H�U����el�U�u�K2�l²�gN��X��=�.R
@��2�� 	A$�I5UU��Z4k�Y��ک��к,�r���[[���l�]��Y���W�R��W���5/2���E�j��,ɽdeD�Jf�n^MedQ���(cV�Uc��UUUWv�F�-&�|'/������>;{~ДG��b�9��$�j�����aB�� �H4Y�_��Y�v�m�Q�����Z����,iq���r���LΎ�K#��Ss�0N���,5y��?�tƦYIJ���C���ğ|OH�4*���P�.=q���_���N��c�dG�;gVF
�''��e��Uo|�0�rO�����<��'B�<o�R���A�дc+�n�k��?����1�83���.�嬓*b��>=���,��ŋ&xb���s����:���lN80��C�y�xL�zg����Ԫ���e�[8Ln��"�e��Su�*X���`�ȧ�fSy�wFQ��&[���ʭ��aߜ[��\�u����S��؟ �Yv>�s'K��TtR�Y2{��d���ϧQ��x�z�k,���o�F�x��b���J�dcDo]J��ON>(�'���������8�U��R��_	'��>͠�;,��<O(�iڔ�1}�G�����^p��7uOB��1�C���;b��R�X��f�I��Y�\f��Ōw��`�9T%���xO�)��'yKZG<f����~MF��㙂G�OZ{�?�!�saeKUTQO�R�R\�*G�X�7n�قܪ���dc���^2��n����c�R�/*ŋ"�l�-��D߿H�[�5����"�k0}�hi�hҌv��ڕO��k��_�b+�{�p2v����hL��T<��x���1��>''Ǔs�����'3���.������lKE�Gt�۸xͨ���}�'�ŷ?=U�_c����׽wO*S���*���H��IQ<i�0R,.P�g�?��y4j�{鯡���bx6e�q3��f��V|�ֻ�1Xڕ�UL+�府k7�'�~,Z��䝺����e�a�UVkv���f�=GZrN�l�Y��QS�&�gᣥ�c�WP�mG%GC]�]G�w&��ǟC�rb���tMd��ӿ�s�ʅ���n�����S�3RG�O����С��s������&3���0fgEI6��i�����?�.�k��)�
U!��)Rc�TF���w$S�	�k�