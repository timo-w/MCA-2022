BZh91AY&SY�Q� \_�Ryg����������`  �    �S�i�@ i� 2  ��41�0�L �F��2d��bh�#0�0Mdh8ɓC�� �� �M4i���&MF&�04ѦF�`�$dO&A0F����mM�mS�R�B�1�I��(�D^$��zO�?W�r9���%��ҿ;��W�?/�Er��1���uh�~[w�z�\�߹i8��E��nT�IwPb�I5���MW,2TSz��TmW=#���
,��������9�z�׻����wi���6߆4��x�-iu��L��v����Ml,��QO��X�}���rִ��\j�S��鐼�4絟eՖ4���'B��S'.S��v�~?�mb���m�ڏ�M��2�u^�9�����\	�5۶ַ�t��\ߑ�������O�Q����.��GLvu�'%%+�����3�v�5ڗSuG���م�T�ёyrTU�U2��z���j�K�Z��-S����뵵}+p���V��RRRa)TR�b��;ރ�%&->��9�d]w5h��*�n`_�}9�X�g�VF,X飺�c���u�S�O��UO�b�UZ��������¬�KFm<��6�z�6\��e��r��Z�[����崲�?U�߻v����ZJ��RĺQ��SUR��Y�j�Ɖ�ɬ�t�Jģ%X��[mU������XU괛i������-����h��#�Q���B@01�@p���Z����bD7�v�~.�fy[�\���O���ь��c;�nۍ��UglY;<�N�8͌d�9׺v�o�����41�y�UK��9��	�D�rB���!E"���w���7��9�.ى����׫��_�-V�8=��S�5��tI>6�������p\����+�93��F��ʦ��>�a��F�]㖺%̾xi�E4��e�^TE�\0a|���#��g��9UUL�`o�|�������2x�-����Tw��/c�[(K�.ar���Yii��l��.�OE�Jy�c6����>|�ݎ��7nv2�b�6��78닶WA�����O�b,�z�y���ԪJo1b����;:=���iODM%���c�6ţE���Ii���D�W)R�)�î>i��*8��.����~5W�(�%��7՜�����ˬb�yF�N��s��ws�'��k/]7I�9�^?A�3�|�:���B��@��d��9��I�[��B���:U
�W�K)���>L/��;JZ�9a3fle�h3<�,��7��zS�a���%�T�UE�%*QE%ĸ��ĩ�g4����^/F#���N�$;U��Qm-�b��KZ��J�bȩ�*Kv��6��3V��vrQbќQ-e�a��L�ц��iH^q�Wu�g��R+��֗x��1���P�]�YPn�:���?��8�\[�	��Ror>���f�}�K`Z(�`;'F���kE���=m�yx�]1�a�ϋ�����iNc�ܪNv	#�%D�&��QH�������û6�׾�y����L��a�`șJU2IH�>�K\�,kJ�*����ܦ�����n
��N�}���c�_�UU��f�y�N���BqNl��96��S��eߛ�}a�G8�kGG�u�G��-W�6��kł`�Ä�H��]�Ӕt�(|(��mp�����Q��:��zw8pP�r9E��c�R����:�ƹQRMn��1��Tw6O�O�W��Ɣ��*��ה��<F���w$S�	���